`ifndef VX_TB_DEFINE_VH
`define VX_TB_DEFINE_VH

`define VX_info(ID, message)    `uvm_info(ID, message, UVM_NONE)
`define VX_warning(ID, message) `uvm_warning(ID, message)
`define VX_error(ID, message)   `uvm_error(ID, message)
`define VX_fatal(ID, message)   `uvm_fatal(ID, message)

`endif // VX_TB_DEFINE_VH



