// Copyright © 2019-2023
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

`include "VX_define.vh"

module VX_execute import VX_gpu_pkg::*; #(
    parameter `STRING INSTANCE_ID = "",
    parameter CORE_ID = 0
) (
    `SCOPE_IO_DECL

    input wire              clk,
    input wire              reset,

`ifdef PERF_ENABLE
    input sysmem_perf_t     sysmem_perf,
    input pipeline_perf_t   pipeline_perf,
`endif

    input base_dcrs_t       base_dcrs,

    // Dcache interface
    VX_lsu_mem_if.master    lsu_mem_if [`NUM_LSU_BLOCKS],

    // dispatch interface
    VX_dispatch_if.slave    dispatch_if [NUM_EX_UNITS * `ISSUE_WIDTH],

    // commit interface
    VX_commit_if.master     commit_if [NUM_EX_UNITS * `ISSUE_WIDTH],

    // scheduler interfaces
    VX_sched_csr_if.slave   sched_csr_if,
    VX_branch_ctl_if.master branch_ctl_if [`NUM_ALU_BLOCKS],
    VX_warp_ctl_if.master   warp_ctl_if,

    // commit interface
    VX_commit_csr_if.slave  commit_csr_if
);

`ifdef EXT_F_ENABLE
    VX_fpu_csr_if fpu_csr_if[`NUM_FPU_BLOCKS]();
`endif

    
    localparam alu_dispatch_start_idx = EX_ALU * `ISSUE_WIDTH;
    localparam alu_dispatch_end_idx   = alu_dispatch_start_idx + `ISSUE_WIDTH - 1;
    localparam alu_commit_start_idx   = EX_ALU * `ISSUE_WIDTH;
    localparam alu_commit_end_idx     = alu_commit_start_idx + `ISSUE_WIDTH - 1;
    
    localparam lsu_dispatch_start_idx = EX_LSU * `ISSUE_WIDTH;
    localparam lsu_dispatch_end_idx   = lsu_dispatch_start_idx + `ISSUE_WIDTH - 1;
    localparam lsu_commit_start_idx   = EX_LSU * `ISSUE_WIDTH;
    localparam lsu_commit_end_idx     = lsu_commit_start_idx + `ISSUE_WIDTH - 1;
    
    localparam fpu_dispatch_start_idx = EX_FPU * `ISSUE_WIDTH;
    localparam fpu_dispatch_end_idx   = fpu_dispatch_start_idx + `ISSUE_WIDTH - 1;
    localparam fpu_commit_start_idx   = EX_FPU * `ISSUE_WIDTH;
    localparam fpu_commit_end_idx     = fpu_commit_start_idx + `ISSUE_WIDTH - 1;

    localparam tcu_dispatch_start_idx = EX_TCU * `ISSUE_WIDTH;
    localparam tcu_dispatch_end_idx   = tcu_dispatch_start_idx + `ISSUE_WIDTH - 1;
    localparam tcu_commit_start_idx   = EX_TCU * `ISSUE_WIDTH;
    localparam tcu_commit_end_idx     = tcu_commit_start_idx + `ISSUE_WIDTH - 1;

    localparam sfu_dispatch_start_idx = EX_SFU * `ISSUE_WIDTH;
    localparam sfu_dispatch_end_idx   = sfu_dispatch_start_idx + `ISSUE_WIDTH - 1;
    localparam sfu_commit_start_idx   = EX_SFU * `ISSUE_WIDTH;
    localparam sfu_commit_end_idx     = sfu_commit_start_idx + `ISSUE_WIDTH - 1;

    VX_alu_unit #(
        .INSTANCE_ID (`SFORMATF(("%s-alu", INSTANCE_ID)))
    ) alu_unit (
        .clk            (clk),
        .reset          (reset),
        .dispatch_if    (dispatch_if[alu_dispatch_end_idx : alu_dispatch_start_idx]), 
        .commit_if      (commit_if[alu_commit_end_idx: alu_commit_start_idx]), 
        .branch_ctl_if  (branch_ctl_if)
    );

    `SCOPE_IO_SWITCH (1);

    VX_lsu_unit #(
        .INSTANCE_ID (`SFORMATF(("%s-lsu", INSTANCE_ID)))
    ) lsu_unit (
        `SCOPE_IO_BIND  (0)
        .clk            (clk),
        .reset          (reset),
        .dispatch_if    (dispatch_if[lsu_dispatch_end_idx : lsu_dispatch_start_idx]),
        .commit_if      (commit_if[lsu_commit_end_idx: lsu_commit_start_idx]), 
        .lsu_mem_if     (lsu_mem_if)
    );

`ifdef EXT_F_ENABLE
    VX_fpu_unit #(
        .INSTANCE_ID (`SFORMATF(("%s-fpu", INSTANCE_ID)))
    ) fpu_unit (
        .clk            (clk),
        .reset          (reset),
        .dispatch_if    (dispatch_if[fpu_dispatch_end_idx : fpu_dispatch_start_idx]), 
        .commit_if      (commit_if[fpu_commit_end_idx : fpu_commit_start_idx]), 
        .fpu_csr_if     (fpu_csr_if)
    );
`endif

`ifdef EXT_TCU_ENABLE
    VX_tcu_unit #(
        .INSTANCE_ID (`SFORMATF(("%s-tcu", INSTANCE_ID)))
    ) tcu_unit (
        .clk            (clk),
        .reset          (reset),
        .dispatch_if    (dispatch_if[tcu_dispatch_end_idx : tcu_dispatch_start_idx]), 
        .commit_if      (commit_if[tcu_commit_end_idx : tcu_commit_start_idx]) 
    );
`endif

    VX_sfu_unit #(
        .INSTANCE_ID (`SFORMATF(("%s-sfu", INSTANCE_ID))),
        .CORE_ID (CORE_ID)
    ) sfu_unit (
        .clk            (clk),
        .reset          (reset),
    `ifdef PERF_ENABLE
        .sysmem_perf    (sysmem_perf),
        .pipeline_perf  (pipeline_perf),
    `endif
        .base_dcrs      (base_dcrs),
        .dispatch_if    (dispatch_if[sfu_dispatch_end_idx : sfu_dispatch_start_idx]), 
        .commit_if      (commit_if[sfu_commit_end_idx : sfu_commit_start_idx]), 
    `ifdef EXT_F_ENABLE
        .fpu_csr_if     (fpu_csr_if),
    `endif
        .commit_csr_if  (commit_csr_if),
        .sched_csr_if   (sched_csr_if),
        .warp_ctl_if    (warp_ctl_if)
    );

endmodule
