class VX_risc_v_seq_item extends uvm_sequence_item;

    rand risc_v_data_type_t           data_type;
    rand risc_v_seq_data_t            raw_data;

    `uvm_object_utils_begin(VX_risc_v_seq_item);    
        `uvm_field_enum(risc_v_data_type_t, data_type,      UVM_ALL_ON)
        `uvm_field_int(raw_data,                            UVM_ALL_ON)
    
    `uvm_object_utils_end

    function new(string name="VX_risc_v_seq_item");
        super.new(name);
    endfunction
  
endclass

class VX_risc_v_inst_seq_item extends VX_risc_v_seq_item;

    rand risc_v_seq_inst_type_t       inst_type;
    rand risc_v_seq_opcode_t          opcode;
    
    `uvm_object_utils_begin(VX_risc_v_inst_seq_item);    
        `uvm_field_enum(risc_v_seq_inst_type_t, inst_type, UVM_ALL_ON)  
        `uvm_field_int(opcode,                             UVM_ALL_ON)
    `uvm_object_utils_end

    function new(string name="VX_risc_v_inst_seq_item");
        super.new(name);
    endfunction
  
endclass

