`ifndef VX_TB_COMMON_PKG_VH
`define VX_TB_COMMON_PKG_VH

package VX_tb_common_pkg;


    `include "VX_tb_types.svh"
    `include "VX_sequence_items.sv"
    
endpackage

`endif // VX_TB_COMMON_PKG_VH
