class VX_execute_tb_txn_item extends uvm_transaction;

    `uvm_object_utils(VX_execute_tb_txn_item)

    function new(string name="VX_execute_tb_txn_item");
        super.new(name);
    endfunction

endclass