`timescale 1ns/1ps

import uvm_pkg::*;
import VX_gpu_pkg::*;